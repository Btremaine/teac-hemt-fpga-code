//////////////////////////////////////////////////////////////////////////////
// Module     : defines.v                                                   //
// Description: This module contains system level definitions.              //
//////////////////////////////////////////////////////////////////////////////

`define NUM_DACS               5'd20
`undef BENCH
//`define BENCH
